module control(
	input logic Reset,
	input logic Clk,
	input logic Run,
	input logic ClearA_LoadB,
	output logic Clr_Ld,
	output logic Shift,
	output logic Add,
	output logic Sub
);


endmodule