module testbench();

timeunit 10ns;	// Half clock cycle at 50 MHz
			// This is the amount of time represented by #1 
timeprecision 1ns;


logic[7:0] Switches;
logic Reset, Run, ClearA_LoadB, X;
logic Clk = 0;

logic[6:0] AhexU;
logic[6:0] AhexL;
logic[6:0] BhexU;
logic[6:0] BhexL;
logic[7:0] Aval;
logic[7:0] Bval;

multiplier_toplevel testee(.S(Switches), .*);

// Toggle the clock
// #1 means wait for a delay of 1 timeunit
always begin: CLOCK_GENERATION
#1 Clk = ~Clk;
end

initial begin: CLOCK_INITIALIZATION
    Clk = 0;
end 

initial begin: testing
	Reset = 1;
	Run = 0;
	ClearA_LoadB = 0;
	
	#2
	Reset = 0;
	#2
	Switches = -8'd5;
	ClearA_LoadB = 1;
	#2
	ClearA_LoadB = 0;
	#4
	Switches = 8'd3;
	#2
	Run = 1;
	#40
	Run = 0;
	#10
	Run = 1;
	#3
	Run = 0;
end

endmodule