module testbench();

timeunit 10ns;	// Half clock cycle at 50 MHz
			// This is the amount of time represented by #1 
timeprecision 1ns;

logic Clk = 0;

// Toggle the clock
// #1 means wait for a delay of 1 timeunit
always begin : CLOCK_GENERATION
#1 Clk = ~Clk;
end

initial begin: CLOCK_INITIALIZATION
    Clk = 0;
end

logic [15:0] S;
logic Reset, Run, Continue;
logic [11:0] LED;
logic [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7;
logic CE, UB, LB, OE, WE;
logic [19:0] ADDR;
wire [15:0] Data;

lab6_toplevel tested(.*);


initial begin : testLoop
	S = 20; //XOR test
	Continue = 0;
	#20 Reset = 1;
	#2 Reset = 0;
	#2 Reset = 1;
	#20 Run = 1;
	#2 Run = 0;
	#2 Run = 1;
	
	//XOR test, expected result is 1010 0101 1010 0101, or A5A5
	#100 S = 16'b1111000011110000;
	Continue = 1;
	#100 S = 16'b0101010101010101;
	Continue = 0;
	#10 Continue = 1;
end

endmodule