module SRAM_controller(
	input logic SRAM_CLK
);

endmodule